magic
tech sky130B
magscale 1 2
timestamp 1762372176
<< nwell >>
rect 752 -654 1272 -560
rect 752 -754 834 -654
rect 868 -754 1272 -654
rect 752 -760 1272 -754
rect 752 -776 912 -760
rect 752 -788 818 -776
rect 752 -834 912 -788
rect 1120 -834 1272 -760
rect 752 -902 1272 -834
rect 752 -904 956 -902
rect 752 -920 852 -904
rect 934 -920 956 -904
rect 754 -1084 816 -1034
rect 990 -1168 1032 -902
rect 1066 -920 1272 -902
rect 754 -1204 790 -1202
rect 990 -1204 1034 -1168
<< ndiff >>
rect 990 -1396 1036 -1392
rect 516 -1464 716 -1424
rect 958 -1536 1066 -1396
rect 1296 -1418 1530 -1398
rect 1296 -1488 1542 -1418
rect 956 -1592 1066 -1536
<< pdiff >>
rect 792 -1084 816 -1034
rect 990 -1168 1032 -964
rect 990 -1204 1034 -1168
<< poly >>
rect 398 -1118 448 -1016
rect 398 -1396 458 -1330
rect 896 -1362 962 -1304
rect 1060 -1354 1126 -1304
rect 1084 -1362 1122 -1360
rect 1576 -1392 1626 -1326
rect 754 -1558 804 -1492
rect 1200 -1558 1250 -1492
rect 802 -1752 852 -1686
<< locali >>
rect 532 -618 1488 -546
rect 532 -1010 696 -618
rect 916 -622 1488 -618
rect 818 -756 874 -654
rect 912 -834 1120 -760
rect 984 -1000 1040 -834
rect 398 -1118 448 -1016
rect 486 -1302 688 -1162
rect 754 -1168 832 -1002
rect 990 -1168 1032 -1000
rect 754 -1206 826 -1168
rect 990 -1204 1034 -1168
rect 508 -1328 666 -1302
rect 398 -1396 448 -1330
rect 754 -1388 792 -1206
rect 896 -1354 962 -1304
rect 1060 -1354 1126 -1304
rect 1214 -1388 1250 -960
rect 1324 -1010 1488 -622
rect 1360 -1162 1512 -1130
rect 1336 -1302 1538 -1162
rect 482 -1424 520 -1416
rect 482 -1438 716 -1424
rect 408 -1464 716 -1438
rect 408 -1498 586 -1464
rect 408 -1650 466 -1498
rect 754 -1596 902 -1388
rect 956 -1396 958 -1392
rect 990 -1396 1036 -1392
rect 1052 -1396 1056 -1392
rect 956 -1598 1066 -1396
rect 1116 -1596 1250 -1388
rect 1576 -1392 1626 -1326
rect 1296 -1418 1530 -1398
rect 1296 -1428 1542 -1418
rect 1296 -1488 1590 -1428
rect 1488 -1498 1590 -1488
rect 408 -1808 690 -1650
rect 802 -1752 852 -1686
rect 970 -1692 1038 -1598
rect 1532 -1658 1590 -1498
rect 886 -1808 1094 -1746
rect 1308 -1808 1590 -1658
rect 408 -1818 1590 -1808
rect 408 -1856 902 -1818
rect 1078 -1856 1590 -1818
rect 408 -1870 1590 -1856
<< viali >>
rect 902 -1856 1078 -1818
<< metal1 >>
rect 820 -660 884 -654
rect 820 -748 826 -660
rect 878 -748 884 -660
rect 820 -754 884 -748
rect 912 -782 1120 -760
rect 912 -834 946 -782
rect 1088 -834 1120 -782
rect 288 -904 358 -898
rect 288 -968 298 -904
rect 350 -968 358 -904
rect 846 -910 942 -904
rect 846 -962 852 -910
rect 936 -962 942 -910
rect 846 -968 942 -962
rect 1080 -908 1176 -902
rect 1080 -960 1086 -908
rect 1170 -960 1176 -908
rect 288 -974 358 -968
rect 288 -1678 354 -974
rect 398 -1116 448 -1016
rect 792 -1084 816 -1034
rect 390 -1122 456 -1116
rect 390 -1186 396 -1122
rect 450 -1186 456 -1122
rect 390 -1192 456 -1186
rect 398 -1330 448 -1192
rect 498 -1276 676 -1162
rect 790 -1204 826 -1144
rect 990 -1168 1032 -964
rect 1080 -966 1176 -960
rect 1188 -1082 1250 -1034
rect 1360 -1162 1366 -1130
rect 990 -1204 1034 -1168
rect 1336 -1180 1366 -1162
rect 1506 -1162 1512 -1130
rect 1506 -1180 1538 -1162
rect 792 -1206 826 -1204
rect 498 -1328 516 -1276
rect 658 -1328 676 -1276
rect 1336 -1302 1538 -1180
rect 1574 -1264 1624 -1016
rect 1566 -1270 1632 -1264
rect 1194 -1304 1246 -1302
rect 398 -1396 458 -1330
rect 498 -1336 676 -1328
rect 776 -1354 962 -1304
rect 776 -1366 828 -1354
rect 896 -1362 962 -1354
rect 1060 -1354 1246 -1304
rect 1566 -1334 1572 -1270
rect 1626 -1334 1632 -1270
rect 1566 -1340 1632 -1334
rect 1060 -1360 1084 -1354
rect 1060 -1362 1122 -1360
rect 764 -1372 828 -1366
rect 600 -1424 620 -1398
rect 486 -1438 716 -1424
rect 408 -1464 716 -1438
rect 764 -1436 770 -1372
rect 822 -1436 828 -1372
rect 1188 -1368 1246 -1354
rect 1188 -1374 1252 -1368
rect 764 -1442 828 -1436
rect 956 -1396 958 -1392
rect 990 -1396 1036 -1392
rect 1052 -1396 1056 -1392
rect 408 -1498 586 -1464
rect 628 -1492 648 -1464
rect 408 -1650 466 -1498
rect 516 -1554 716 -1552
rect 516 -1606 524 -1554
rect 700 -1606 716 -1554
rect 754 -1558 804 -1492
rect 956 -1592 1066 -1396
rect 1188 -1438 1194 -1374
rect 1246 -1438 1252 -1374
rect 1574 -1392 1626 -1340
rect 1188 -1444 1252 -1438
rect 1296 -1418 1530 -1398
rect 1296 -1428 1542 -1418
rect 1296 -1488 1590 -1428
rect 1200 -1558 1250 -1492
rect 1488 -1498 1590 -1488
rect 1296 -1550 1484 -1544
rect 516 -1612 716 -1606
rect 1296 -1602 1302 -1550
rect 1478 -1602 1484 -1550
rect 1296 -1608 1484 -1602
rect 288 -1688 358 -1678
rect 288 -1752 298 -1688
rect 350 -1752 358 -1688
rect 288 -1758 358 -1752
rect 408 -1808 690 -1650
rect 1532 -1658 1590 -1498
rect 790 -1686 850 -1680
rect 844 -1752 852 -1686
rect 790 -1758 850 -1752
rect 890 -1808 1090 -1782
rect 1308 -1808 1590 -1658
rect 408 -1818 1590 -1808
rect 408 -1856 902 -1818
rect 1078 -1856 1590 -1818
rect 408 -1870 1590 -1856
<< via1 >>
rect 826 -748 878 -660
rect 946 -834 1088 -782
rect 298 -968 350 -904
rect 852 -962 936 -910
rect 1086 -960 1170 -908
rect 396 -1186 450 -1122
rect 1366 -1180 1506 -1128
rect 516 -1328 658 -1276
rect 1572 -1334 1626 -1270
rect 770 -1436 822 -1372
rect 524 -1606 700 -1554
rect 1194 -1438 1246 -1374
rect 1302 -1602 1478 -1550
rect 298 -1752 350 -1688
rect 790 -1752 844 -1686
<< metal2 >>
rect 474 -660 884 -654
rect 474 -748 826 -660
rect 878 -748 884 -660
rect 474 -754 884 -748
rect 912 -782 1098 -776
rect 912 -788 946 -782
rect 480 -834 946 -788
rect 1088 -834 1098 -782
rect 480 -840 1098 -834
rect 288 -902 358 -898
rect 288 -904 1176 -902
rect 288 -968 298 -904
rect 350 -908 1176 -904
rect 350 -910 1086 -908
rect 350 -962 852 -910
rect 936 -960 1086 -910
rect 1170 -960 1176 -908
rect 936 -962 1176 -960
rect 350 -966 1176 -962
rect 350 -968 1080 -966
rect 288 -974 358 -968
rect 390 -1122 456 -1116
rect 1336 -1122 1528 -1118
rect 390 -1186 396 -1122
rect 450 -1126 1528 -1122
rect 450 -1182 1342 -1126
rect 1518 -1182 1528 -1126
rect 450 -1186 1528 -1182
rect 390 -1192 456 -1186
rect 1336 -1192 1528 -1186
rect 506 -1270 666 -1262
rect 1566 -1270 1632 -1264
rect 506 -1272 1572 -1270
rect 506 -1328 516 -1272
rect 658 -1328 1572 -1272
rect 506 -1334 1572 -1328
rect 1626 -1334 1632 -1270
rect 506 -1336 1632 -1334
rect 506 -1338 666 -1336
rect 1566 -1340 1632 -1336
rect 764 -1372 828 -1366
rect 764 -1374 770 -1372
rect 346 -1428 770 -1374
rect 764 -1436 770 -1428
rect 822 -1436 828 -1372
rect 764 -1442 828 -1436
rect 1188 -1374 1252 -1368
rect 1188 -1438 1194 -1374
rect 1246 -1384 1252 -1374
rect 1246 -1438 1694 -1384
rect 1188 -1444 1252 -1438
rect 514 -1552 710 -1544
rect 1292 -1546 1488 -1536
rect 514 -1608 524 -1552
rect 700 -1608 712 -1552
rect 514 -1612 712 -1608
rect 1292 -1602 1300 -1546
rect 1476 -1550 1488 -1546
rect 1478 -1602 1488 -1550
rect 1292 -1612 1488 -1602
rect 514 -1618 710 -1612
rect 288 -1680 358 -1678
rect 288 -1686 850 -1680
rect 288 -1688 790 -1686
rect 288 -1752 298 -1688
rect 350 -1752 790 -1688
rect 844 -1752 850 -1686
rect 288 -1758 850 -1752
<< via2 >>
rect 1342 -1128 1518 -1126
rect 1342 -1180 1366 -1128
rect 1366 -1180 1506 -1128
rect 1506 -1180 1518 -1128
rect 1342 -1182 1518 -1180
rect 516 -1276 658 -1272
rect 516 -1328 658 -1276
rect 524 -1554 700 -1552
rect 524 -1606 700 -1554
rect 524 -1608 700 -1606
rect 1300 -1550 1476 -1546
rect 1300 -1602 1302 -1550
rect 1302 -1602 1476 -1550
<< metal3 >>
rect 1336 -1126 1528 -1118
rect 1336 -1182 1342 -1126
rect 1518 -1182 1528 -1126
rect 1336 -1192 1528 -1182
rect 506 -1272 666 -1262
rect 506 -1328 516 -1272
rect 658 -1328 666 -1272
rect 506 -1338 666 -1328
rect 524 -1544 658 -1338
rect 1342 -1536 1488 -1192
rect 514 -1552 710 -1544
rect 514 -1608 524 -1552
rect 700 -1608 710 -1552
rect 514 -1618 710 -1608
rect 1292 -1546 1488 -1536
rect 1292 -1602 1300 -1546
rect 1476 -1602 1488 -1546
rect 1292 -1612 1488 -1602
use sky130_fd_pr__nfet_01v8_9ZWGZ9  sky130_fd_pr__nfet_01v8_9ZWGZ9_0
timestamp 1760634725
transform -1 0 1093 0 1 -1461
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_9ZWGZ9  sky130_fd_pr__nfet_01v8_9ZWGZ9_1
timestamp 1760634725
transform 0 -1 959 1 0 -1719
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_9ZWGZ9  sky130_fd_pr__nfet_01v8_9ZWGZ9_2
timestamp 1760634725
transform -1 0 929 0 1 -1461
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_9ZWGZ9  sky130_fd_pr__nfet_01v8_9ZWGZ9_3
timestamp 1760634725
transform 0 1 647 -1 0 -1525
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_ML4XRG  sky130_fd_pr__nfet_01v8_ML4XRG_0
timestamp 1761100160
transform 0 1 555 -1 0 -1363
box -73 -157 73 157
use sky130_fd_pr__nfet_01v8_ML4XRG  sky130_fd_pr__nfet_01v8_ML4XRG_1
timestamp 1761100160
transform 0 -1 1469 1 0 -1361
box -73 -157 73 157
use sky130_fd_pr__pfet_01v8_KDZMJM  sky130_fd_pr__pfet_01v8_KDZMJM_0
timestamp 1761100160
transform 0 1 1470 -1 0 -1066
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_KDZMJM  sky130_fd_pr__pfet_01v8_KDZMJM_1
timestamp 1761100160
transform 1 0 1128 0 1 -1066
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_KDZMJM  sky130_fd_pr__pfet_01v8_KDZMJM_2
timestamp 1761100160
transform 0 -1 552 1 0 -1066
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_KDZMJM  sky130_fd_pr__pfet_01v8_KDZMJM_3
timestamp 1761100160
transform 0 -1 982 1 0 -706
box -144 -198 144 164
use sky130_fd_pr__pfet_01v8_KDZMJM  XMmirr3
timestamp 1761100160
transform 1 0 894 0 1 -1066
box -144 -198 144 164
use sky130_fd_pr__nfet_01v8_9ZWGZ9  Xsky130_fd_pr__nfet_01v8_9ZWGZ9_1
timestamp 1760634725
transform 0 -1 1357 1 0 -1525
box -73 -157 73 157
<< labels >>
rlabel metal2 346 -1428 770 -1374 1 Vm
rlabel metal2 1246 -1438 1694 -1384 1 vp
rlabel metal2 480 -840 946 -788 1 vdd
rlabel metal2 474 -754 826 -654 1 vbias_p
rlabel metal2 658 -1336 1572 -1270 1 voutp
rlabel metal2 450 -1186 1366 -1122 1 voutn
flabel metal1 886 -1870 1086 -1842 0 FreeSans 80 0 0 0 gnd
port 3 nsew
rlabel metal2 288 -1758 358 -1678 1 vbias_n
<< end >>
