** sch_path: /home/user/projects/nic2025_v2/nic2025_openDVS/analog/xschem/final/col_amp_n_clamp_v1/col_amp_v1.sch
**.subckt col_amp_v1 vdd pbias pbchk vcascp vout_sense pix_rst vcascn gnd bias_amp_cascn feedback sense
*.iopin vdd
*.iopin gnd
*.iopin sense
*.iopin vout_sense
*.iopin feedback
*.iopin pbchk
*.iopin pix_rst
*.iopin vcascn
*.iopin vcascp
*.iopin pbias
*.iopin bias_amp_cascn
XMpb pbchk pbias vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 ad=1.45 as=1.45 pd=10.58 ps=10.58 nrd=0.058 nrs=0.058 sa=0 sb=0 sd=0
+ mult=1 m=1
XMnc vout_sense amp_p_vg sense gnd sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 ad=0.87 as=0.87 pd=6.58 ps=6.58 nrd=0.0966666666666667
+ nrs=0.0966666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XMfb vout_sense pix_rst feedback gnd sky130_fd_pr__nfet_01v8 L=0.5 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58
+ sa=0 sb=0 sd=0 mult=1 m=1
XMpc vout_sense vcascp pbchk vdd sky130_fd_pr__pfet_01v8 L=1 W=5 nf=1 ad=1.45 as=1.45 pd=10.58 ps=10.58 nrd=0.058 nrs=0.058 sa=0
+ sb=0 sd=0 mult=1 m=1
x1 vdd amp_p_vg vcascn sense bias_amp_cascn gnd amp_p_5T
**.ends

* expanding   symbol:  /home/user/projects/open_dvs/analog/amp_p_5T.sym # of pins=6
** sym_path: /home/user/projects/open_dvs/analog/amp_p_5T.sym
** sch_path: /home/user/projects/open_dvs/analog/amp_p_5T.sch
.subckt amp_p_5T vdd vout vp vm vbias gnd
*.iopin gnd
*.iopin vdd
*.iopin vout
*.iopin vm
*.iopin vp
*.iopin vbias
XMinm vout vm vsource vdd sky130_fd_pr__pfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMinp vdio vp vsource vdd sky130_fd_pr__pfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMdio vdio vdio gnd gnd sky130_fd_pr__nfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMmirr vout vdio gnd gnd sky130_fd_pr__nfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMbias vsource vbias vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
.ends

.end
