** sch_path: /home/user/projects/nic2025_v2/nic2025_openDVS/analog/xschem/final/col_amp_n_clamp_v1/clamp_qdvs_v2.sch
**.subckt clamp_qdvs_v2 vdd clamp_leakp CLAMP_RST vgn vout vamp vcm vgp _CLAMP_RST clamp_leakn gnd
*.iopin vdd
*.iopin gnd
*.iopin vcm
*.iopin _CLAMP_RST
*.iopin CLAMP_RST
*.iopin clamp_leakp
*.iopin clamp_leakn
*.iopin vout
*.iopin vamp
*.opin vgn
*.opin vgp
XM1 vgn vgn vcm gnd sky130_fd_pr__nfet_01v8 L=0.5 W=0.75 nf=1 ad=0.2175 as=0.2175 pd=2.08 ps=2.08 nrd=0.386666666666667
+ nrs=0.386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM2 vgp vgp vcm vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM3 vgn clamp_leakp vdd vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM4 vgp clamp_leakn gnd gnd sky130_fd_pr__nfet_01v8 L=0.5 W=0.75 nf=1 ad=0.2175 as=0.2175 pd=2.08 ps=2.08 nrd=0.386666666666667
+ nrs=0.386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM5 vdd vgn vout gnd sky130_fd_pr__nfet_01v8 L=0.5 W=0.75 nf=1 ad=0.2175 as=0.2175 pd=2.08 ps=2.08 nrd=0.386666666666667
+ nrs=0.386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM6 gnd vgp vout vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
XM7 vout _CLAMP_RST vamp gnd sky130_fd_pr__nfet_01v8 L=0.5 W=0.75 nf=1 ad=0.2175 as=0.2175 pd=2.08 ps=2.08 nrd=0.386666666666667
+ nrs=0.386666666666667 sa=0 sb=0 sd=0 mult=1 m=1
XM8 vout CLAMP_RST vamp vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1.5 nf=1 ad=0.435 as=0.435 pd=3.58 ps=3.58 nrd=0.193333333333333
+ nrs=0.193333333333333 sa=0 sb=0 sd=0 mult=1 m=1
**.ends
.end
