** sch_path: /home/user/projects/nic2025_v2/nic2025_openDVS/analog/xschem/final/col_amp_n_clamp_v1/amp_p_5T.sch
**.subckt amp_p_5T vdd vout vp vm vbias gnd
*.iopin gnd
*.iopin vdd
*.iopin vout
*.iopin vm
*.iopin vp
*.iopin vbias
XMinm vout vm vsource vdd sky130_fd_pr__pfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMinp vdio vp vsource vdd sky130_fd_pr__pfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMdio vdio vdio gnd gnd sky130_fd_pr__nfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMmirr vout vdio gnd gnd sky130_fd_pr__nfet_01v8 L=0.2 W=0.5 nf=1 ad=0.145 as=0.145 pd=1.58 ps=1.58 nrd=0.58 nrs=0.58 sa=0 sb=0
+ sd=0 mult=1 m=1
XMbias vsource vbias vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
**.ends
.end
